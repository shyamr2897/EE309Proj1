library ieee;
use ieee.std_logic_1164.all;
package mem_package is
type arr is array (65535 downto 0) of std_logic_vector(7 downto 0);
constant MEM_INIT : arr:= (
0 => "10101011",
1 => "00110010",
2 => "01010100",
3 => "00110101",
4 => "01011000",
5 => "00000100",
6 => "11001001",
7 => "00100100",
8 => "00000010",
9 => "00010111",
10 => "01011010",
11 => "00000100",
12 => "00101000",
13 => "00100111",
14 => "11111111",
15 => "00111101",
16 => "10101000",
17 => "00101011",
18 => "00001001",
19 => "00000111",
20 => "11010010",
21 => "00101010",
22 => "11000010",
23 => "11000100",
24 => "00000010",
25 => "00111110",
26 => "11111111",
27 => "00111100",
28 => "11111111",
29 => "00111000",
30 => "00001001",
31 => "00101101",
others => (others => '0'));
end package mem_package;
